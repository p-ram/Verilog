module top_module( output one, output zero );

// Insert your code here
    assign one = 1;
    assign zero=0;

endmodule
