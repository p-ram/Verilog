module top_module(input in, output out);
  
  //wire in verilog is directional, below statement is contineous assignment
  assign out=in;
  
endmodule
